library ieee;
use ieee.std_logic_1164.all;

entity single_cycle is
	generic
	(
	
	);
	port
	(
	
	);
end single_cycle;


architecture Structure of single_cycle is 
	component 
	generic
	(
	
	);
	port
	(
	
	);
	end component;
begin
	
end Structure;